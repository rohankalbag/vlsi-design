CMOS Inverter Transfer Characteristics

.include models-180nm

*Name: Rohan Rajesh Kalbag 
*Roll 20D170033 :  nn = 33

*geometry parameters
.param pw = 1.505U
.param pl = 0.18U
.param pad = {2*pw*pl}
.param pas = {2*pw*pl}
.param ppd = {2*(pw + 2*pl)}
.param pps = {2*(pw + 2*pl)}

.param nw = 0.502U
.param nl = 0.18U
.param nad = {2*nw*nl}
.param nas = {2*nw*nl}
.param npd = {2*(nw + 2*nl)}
.param nps = {2*(nw + 2*nl)}

* unit inverter
.subckt inv supply Inp Output
MP1 Output Inp Supply Supply cmosp
+ L={pl} W={pw} AD={pad} AS={pas} PD={ppd} PS={pps}
MN1 Output Inp 0 0 cmosn
+ L={nl} W={nw} AD={nad} AS={nas} PD={npd} PS={nps}
.ends

vdd supply 0 dc 1.8
* device under test
x3 supply Ck dutout inv
* load capacitor
C3 dutout 0 0.05pF
*transient analysis with pulse inputs
VCk Ck 0 DC

.dc VCk 0 1.8 0.001
.control
run

*plotting of graphs
plot V(dutout) vs V(Ck)
plot deriv(V(dutout)) vs V(Ck)

*calculation of noise margin
let der = deriv(V(dutout))
meas dc VIL find V(Ck) when der = -1
meas dc VIH find V(Ck) when der = -1 rise = last
meas dc VOH find V(dutout) when V(ck) = VIL
meas dc VOL find V(dutout) when V(ck) = VIH

let highnoisemargin = VOH - VIH
let lownoisemargin = VIL - VOL

print highnoisemargin
print lownoisemargin
.endc
.end