Assignment 3

.include models-180nm

*Name: Rohan Rajesh Kalbag 
*Roll 20D170033 :  nn = 33

*geometry parameters
.param pw = 1.505U
.param pl = 0.18U
.param pad = {2*pw*pl}
.param pas = {2*pw*pl}
.param ppd = {2*(pw + 2*pl)}
.param pps = {2*(pw + 2*pl)}

.param nw = 0.502U
.param nl = 0.18U
.param nad = {2*nw*nl}
.param nas = {2*nw*nl}
.param npd = {2*(nw + 2*nl)}
.param nps = {2*(nw + 2*nl)}

* unit inverter from assignment 1 
.subckt inv supply Inp Output
MP1 Output Inp Supply Supply cmosp
+ L={pl} W={pw} AD={pad} AS={pas} PD={ppd} PS={pps}
MN1 Output Inp 0 0 cmosn
+ L={nl} W={nw} AD={nad} AS={nas} PD={npd} PS={nps}
.ends

* pulse with time period of Trep, rise and fall times = Trep/20
.param Trep= 5n
.param Trf = {Trep/20.0}
.param Tw = {Trep/2.0 - Trf}
.param hival=1.8
.param loval=0.0
Vpulse pgen 0 DC 0 PULSE({loval} {hival} {Tw} {Trf} {Trf} {Tw} {Trep})

vdd supply 0 dc 1.8
x1 supply pgen n1 inv
x2 supply n1 n2 inv
x3 supply n2 dutin inv

*input shapers
xi1 supply n2 n3 inv
xi2 supply n2 n3 inv
xi3 supply n2 n3 inv
c1 n3 0 0.1p

*dut 
xdut supply dutin dutout inv

*test load
xl1 supply dutout n4 inv
xl2 supply dutout n4 inv
xl3 supply dutout n4 inv
xl4 supply dutout n4 inv
xl5 supply dutout n4 inv
xl6 supply dutout n4 inv
xl7 supply dutout n4 inv
xl8 supply dutout n4 inv

*load on load 
xll1 supply n4 n5 inv
xll2 supply n4 n5 inv
xll3 supply n4 n5 inv
xll4 supply n4 n5 inv
c2 n5 0 0.1p

.tran 0.1pS {3*Trep} 0nS
.control

run
plot v(dutin) v(dutout)
meas tran delay_rising_edge TRIG v(dutin) VAL=0.9 RISE=2 TARG v(dutout) VAL=0.9 FALL=2
meas tran delay_falling_edge TRIG v(dutin) VAL=0.9 FALL=2 TARG v(dutout) VAL=0.9 RISE=2
let delay = {(delay_rising_edge + delay_falling_edge)/2}
print delay

let gamma = {1.505u/0.502u}
print gamma
.endc
.end